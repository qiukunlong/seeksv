@left_chr	left_pos	left_strand	left_clip_read_NO	right_chr	right_pos	right_strand	right_clip_read_NO	microhomology_length	abnormal_readpair_NO	svtype	left_pos_depth	right_pos_depth	average_depth_of_left_pos_5end	average_depth_of_left_pos_3end	average_depth_of_right_pos_5end	average_depth_of_right_pos_3end	left_pos_clip_percentage	right_pos_clip_percentage	left_seq_cigar	right_seq_cigar	left_seq	right_seq	left_clip_read_NO_of_control	right_clip_read_NO_of_control	abnormal_read_pair_no_of_control
chr17	495	+	17	chr17	700	+	18	4	52	DEL	35	29	15	0	0	27	1	1.2069	79M	4S42M	CATAAATAATACTGGTTTATTACAGAAGCACTAGAAAATGCATGTGGACAAAAGTTGGGATTAGGAGAAAGAAATGAAG	GCATAAAGAAGCCGGACTCACAGGGCAACACACTATCTGACTGTTT	0	0	0
