@left_chr	left_pos	left_strand	left_clip_read_NO	right_chr	right_pos	right_strand	right_clip_read_NO	microhomology_length	abnormal_readpair_NO	svtype	left_pos_depth	right_pos_depth	average_depth_of_left_pos_5end	average_depth_of_left_pos_3end	average_depth_of_right_pos_5end	average_depth_of_right_pos_3end	left_pos_clip_percentage	right_pos_clip_percentage	left_seq_cigar	right_seq_cigar	left_seq	right_seq
chr17	495	+	17	chr17	700	+	18	4	52	DEL	35	29	15	0	0	27	1	1.2069	79M	4S42M	CATAAATAATACTGGTTTATTACAGAAGCACTAGAAAATGCATGTGGACAAAAGTTGGGATTAGGAGAAAGAAATGAAG	GCATAAAGAAGCCGGACTCACAGGGCAACACACTATCTGACTGTTT
chr17	1950	+	18	chr17	2251	+	15	0	54	DEL	29	27	27	0	0	26	1.13793	1.22222	66M	97M	CCGCCCTGTGCCGTGTACCTCTGAGCCCTCTGCACAGTGCCTTCTGCTTGCCTGTGGCTTTGAGAA	AGATGAGCTTTATAAAAATAATGGTGCTAGCTGGGCATGGTGGCTTGCACCTGTAATCCCAGCACTTTGGGAGGCCGAGCTAGGAGGATCGTTTGAG
chr17	4950	+	14	chr17	5151	+	23	0	56	DEL	31	34	28	0	0	29	1.19355	1.08824	68M	97M	AAACTCCTGGGTTCAAGCAATCCTCTCAAGTAGTTAGGACTACAGGGACATGCCACTACACCAGGCTA	CACGAGGAGTACTGGCCTCTTCATGGTGCCAAGATGTCCCTGAGGCCTTAGTCACCTGGGTCCTTGGTGTCCCCTAGGTCAGGGCCATCCCTCTGTC
