@left_chr	left_pos	left_strand	left_clip_read_NO	right_chr	right_pos	right_strand	right_clip_read_NO	microhomology_length	abnormal_readpair_NO	svtype	left_pos_depth	right_pos_depth	average_depth_of_left_pos_5end	average_depth_of_left_pos_3end	average_depth_of_right_pos_5end	average_depth_of_right_pos_3end	left_pos_clip_percentage	right_pos_clip_percentage	left_seq_cigar	right_seq_cigar	left_seq	right_seq
chr17	1950	+	20	chr17	2251	+	28	0	60	DEL	43	43	32	0	0	31	1.11628	1.11628	69M	94M	GAGCCGCCCTGTGCCGTGTACCTCTGAGCCCTCTGCACAGTGCCTTCTGCTTGCCTGTGGCTTTGAGAA	AGATGAGCTTTATAAAAATAATGGTGCTAGCTGGGCATGGTGGCTTGCACCTGTAATCCCAGCACTTTGGGAGGCCGAGCTAGGAGGATCGTTT
chr17	4950	+	17	chr17	5151	+	17	0	50	DEL	28	30	28	0	0	27	1.21429	1.13333	68M	97M	AAATTCCTGGGTGCAAGCAATCCTCTCAAGTAGTTAGGACTACAGGGACATGCCACTACACCAGGCTA	CACGAGGAGTACTGGCCTCTTCATGGTGCCAAGATGTCCCTGAGGCCTTAGTCACCTGGGTCCTTGGTGTCCCCTAGGTCAGGGCCATCCCTCTGTC
